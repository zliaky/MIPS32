`include "defines.v"
module openmips(
	input		wire					clk,
	input		wire					rst,

	input		wire[5:0]				int_i,

	//wishbone����
	input		wire[`RegBus]			wishbone_data_i,
	input		wire					wishbone_ack_i,
	output		wire[`RegBus]			wishbone_addr_o,
	output		wire[`RegBus]			wishbone_data_o,
	output		wire					wishbone_we_o,
	output		wire[15:0]				wishbone_select_o,

	output		wire					timer_int_o,

	input		wire[31:0]				select,
	output		wire[31:0]				data_o
	);

	//����IF/IDģ��������׶�IDģ��ı���
	wire[`InstAddrBus]		pc;
	wire[`InstBus]			inst_i;
	wire[`InstAddrBus]		id_pc_i;
	wire[`InstBus]			id_inst_i;
	wire[`InstAddrBus]		next_pc;

	//��������׶�IDģ�������ID/EXģ�������ı���
	wire[`AluOpBus]			id_aluop_o;
	wire[`AluSelBus]		id_alusel_o;
	wire[`RegBus]			id_reg1_o;
	wire[`RegBus]			id_reg2_o;
	wire					id_wreg_o;
	wire[`RegAddrBus]		id_wd_o;
	wire					id_is_in_delayslot_o;
	wire[`RegBus]			id_link_address_o;
	wire[`RegBus]			id_inst_o;
	wire[31:0]				id_excepttype_o;
	wire[`RegBus]			id_current_inst_address_o;

	//����ID/EXģ�������ִ�н׶�EXģ�������ı���
	wire[`AluOpBus]			ex_aluop_i;
	wire[`AluSelBus]		ex_alusel_i;
	wire[`RegBus]			ex_reg1_i;
	wire[`RegBus]			ex_reg2_i;
	wire					ex_wreg_i;
	wire[`RegAddrBus]		ex_wd_i;
	wire					ex_is_in_delayslot_i;
	wire[`RegBus]			ex_link_address_i;
	wire[`RegBus]			ex_inst_i;
	wire[31:0]				ex_excepttype_i;
	wire[`RegBus]			ex_current_inst_address_i;

	//����ִ�н׶�EX��ģ��������EX/MEMģ�������ı���
	wire					ex_wreg_o;
	wire[`RegAddrBus]		ex_wd_o;
	wire[`RegBus]			ex_wdata_o;
	wire[`RegBus]			ex_hi_o;
	wire[`RegBus]			ex_lo_o;
	wire					ex_whilo_o;
	wire[`AluOpBus]			ex_aluop_o;
	wire[`RegBus]			ex_mem_addr_o;
	wire[`RegBus]			ex_reg1_o;
	wire[`RegBus]			ex_reg2_o;
	wire					ex_cp0_reg_we_o;
	wire[4:0]				ex_cp0_reg_write_addr_o;
	wire[`RegBus]			ex_cp0_reg_data_o;
	wire[31:0]				ex_excepttype_o;
	wire[`RegBus]			ex_current_inst_address_o;
	wire					ex_is_in_delayslot_o;

	//����EX/MEMģ��������ô�׶�MEMģ�������ı���
	wire					mem_wreg_i;
	wire[`RegAddrBus]		mem_wd_i;
	wire[`RegBus]			mem_wdata_i;
	wire[`RegBus]			mem_hi_i;
	wire[`RegBus]			mem_lo_i;
	wire					mem_whilo_i;

	wire[`AluOpBus]			mem_aluop_i;
	wire[`RegBus]			mem_mem_addr_i;
	wire[`RegBus]			mem_reg1_i;
	wire[`RegBus]			mem_reg2_i;	
	wire					mem_cp0_reg_we_i;
	wire[4:0]				mem_cp0_reg_write_addr_i;
	wire[`RegBus] 			mem_cp0_reg_data_i;
	wire[31:0]				mem_excepttype_i;
	wire					mem_is_in_delayslot_i;
	wire[`RegBus]			mem_current_inst_address_i;

	//���ӷô�׶�MEMģ��������MEM/WBģ�������ı���
	wire					mem_wreg_o;
	wire[`RegAddrBus]		mem_wd_o;
	wire[`RegBus]			mem_wdata_o;
	wire[`RegBus]			mem_hi_o;
	wire[`RegBus]			mem_lo_o;
	wire					mem_whilo_o;
	wire 					mem_cp0_reg_we_o;
	wire[4:0] 				mem_cp0_reg_write_addr_o;
	wire[`RegBus] 			mem_cp0_reg_data_o;
	wire[31:0]				mem_excepttype_o;
	wire					mem_is_in_delayslot_o;
	wire[`RegBus]			mem_current_inst_address_o;
	wire[`RegBus]			bad_v_addr_o;

	//����MEM/WBģ���������д�׶ε�����ı���
	wire					wb_wreg_i;
	wire[`RegAddrBus]		wb_wd_i;
	wire[`RegBus]			wb_wdata_i;
	wire[`RegBus]			wb_hi_i;
	wire[`RegBus]			wb_lo_i;
	wire					wb_whilo_i;
	wire 					wb_cp0_reg_we_i;
	wire[4:0] 				wb_cp0_reg_write_addr_i;
	wire[`RegBus] 			wb_cp0_reg_data_i;	
	wire[31:0]				wb_excepttype_i;
	wire					wb_is_in_delayslot_i;
	wire[`RegBus]			wb_current_inst_address_i;

	//��������׶�IDģ����ͨ�üĴ���Regfileģ��ı���
	wire					reg1_read;
	wire					reg2_read;
	wire[`RegBus]			reg1_data;
	wire[`RegBus]			reg2_data;
	wire[`RegAddrBus]		reg1_addr;
	wire[`RegAddrBus]		reg2_addr;

	//����ִ�н׶���hiloģ����������ȡHI��LO�Ĵ���
	wire[`RegBus]			hi;
	wire[`RegBus]			lo;
	
	wire[`DoubleRegBus]		hilo_temp_o;
	wire[1:0]				cnt_o;
	
	wire[`DoubleRegBus]		hilo_temp_i;
	wire[1:0]				cnt_i;
	
	wire					is_in_delayslot_i;
	wire					is_in_delayslot_o;
	wire					next_inst_in_delayslot_o;
	wire					id_branch_flag_o;
	wire[`RegBus]			branch_target_address;
	wire[5:0]				stall;
	wire					stallreq_from_if;
	wire					stallreq_from_id;
	wire					stallreq_from_ex;
	wire					stallreq_from_mem;

	wire[`RegBus]			cp0_data_o;
	wire[4:0]				cp0_raddr_i;

	wire					flush;
	wire[`RegBus]			new_pc;

	wire[`RegBus]			cp0_index;
	wire[`RegBus]			cp0_entry_lo_0;
	wire[`RegBus]			cp0_entry_lo_1;
	wire[`RegBus]			cp0_bad_v_addr;
	wire[`RegBus]			cp0_count;
	wire[`RegBus]			cp0_entry_hi;
	wire[`RegBus]			cp0_compare;
	wire[`RegBus]			cp0_status;
	wire[`RegBus]			cp0_cause;
	wire[`RegBus]			cp0_epc;
	wire[`RegBus]			cp0_ebase;

	wire[`RegBus]			latest_epc;

	wire					rom_ce;

	wire[`RegBus]			ram_addr_o;
	wire					ram_we_o;
	wire[3:0]				ram_sel_o;
	wire[`RegBus]			ram_data_o;
	wire					ram_ce_o;
	wire[`RegBus]			ram_data_i;

	wire[`RegBus]			mmu_addr_i;
	wire[15:0]				mmu_select_i;

	wire[`RegBus]			bus_addr_i;
	wire					bus_write_i;
	wire					tlb_ce_i;
	wire[`RegBus]			tlb_addr_i;

	wire					tlb_we;
	wire[`TLBIndexBus]		tlb_index;
	wire[`TLBDataBus]		tlb_data;
	wire					tlb_excepttype_is_tlbm;
	wire					tlb_excepttype_is_tlbl;
	wire					tlb_excepttype_is_tlbs;

	wire[31:0]				regfile_data_o;
	wire[4:0]				state;
	wire[`InstAddrBus] latch_pc;

	reg[31:0] data_output;
	assign data_o = data_output;
	always @ (*) begin
		if (select[16] == 1'b1) begin
			data_output <= 32'h12345678;
		end else if (select[17] == 1'b1) begin
			data_output <= {31'b0, id_branch_flag_o};
		end else if (select[18] == 1'b1) begin
			data_output <= pc;
		end else if (select[19] == 1'b1) begin
			data_output <= id_inst_i;
		end else if (select[20] == 1'b1) begin
			data_output <= mem_excepttype_o;
		end else if (select[21] == 1'b1) begin
			data_output <= {26'b0, stall};
		end else if (select[22] == 1'b1) begin
			data_output <= {16'b0, mmu_select_i};
		end else if (select[23] == 1'b1) begin
			data_output <= {27'b0, state};
		end else if (select[24] == 1'b1) begin
			data_output <= {31'b0, rst};
		end else if (select[25] == 1'b1) begin
			data_output <= {31'b0, flush};
		end else if (select[26] == 1'b1) begin
			data_output <= next_pc;
		end else if (select[27] == 1'b1) begin
			data_output <= latch_pc;
		end else begin
			data_output <= regfile_data_o;
		end
	end

	//pc_reg����
	pc_reg pc_reg0(
		.clk(clk),
		.rst(rst),
		.stall(stall),
		.flush(flush),
		.new_pc(new_pc),
		.branch_flag_i(id_branch_flag_o),
		.branch_target_address_i(branch_target_address),
		.pc(pc),
		.ce(rom_ce),
		.next_pc(next_pc),
		.latch_pc(latch_pc)
	);

	//IF/IDģ������
	if_id if_id0(
		.clk(clk),
		.rst(rst),
		.stall(stall),
		.flush(flush),
		.if_pc(pc),
		.if_inst(inst_i),
		.id_pc(id_pc_i),
		.id_inst(id_inst_i)
	);

	//����׶�IDģ������
	id id0(
		.rst(rst),
		.pc_i(id_pc_i),
		.inst_i(id_inst_i),
		.ex_aluop_i(ex_aluop_o),

		//����Regfileģ�������
		.reg1_data_i(reg1_data),
		.reg2_data_i(reg2_data),

		//����ִ�н׶ε�ָ��Ҫд���Ŀ�ļĴ�����Ϣ
		.ex_wreg_i(ex_wreg_o),
		.ex_wdata_i(ex_wdata_o),
		.ex_wd_i(ex_wd_o),

		//���ڷô�׶ε�ָ��Ҫд���Ŀ�ļĴ�����Ϣ
		.mem_wreg_i(mem_wreg_o),
		.mem_wdata_i(mem_wdata_o),
		.mem_wd_i(mem_wd_o),

		.is_in_delayslot_i(is_in_delayslot_i),
		//�͵�Regfileģ�����Ϣ
		.reg1_read_o(reg1_read),
		.reg2_read_o(reg2_read),
		.reg1_addr_o(reg1_addr),
		.reg2_addr_o(reg2_addr),

		//�͵�ID/EXģ�����Ϣ
		.aluop_o(id_aluop_o),
		.alusel_o(id_alusel_o),
		.reg1_o(id_reg1_o),
		.reg2_o(id_reg2_o),
		.wd_o(id_wd_o),
		.wreg_o(id_wreg_o),
		.excepttype_o(id_excepttype_o),
		.inst_o(id_inst_o),

		.next_inst_in_delayslot_o(next_inst_in_delayslot_o),
		.branch_flag_o(id_branch_flag_o),
		.branch_target_address_o(branch_target_address),
		.link_addr_o(id_link_address_o),

		.is_in_delayslot_o(id_is_in_delayslot_o),
		.current_inst_address_o(id_current_inst_address_o),
		.stallreq(stallreq_from_id)
	);

	//ͨ�üĴ���Regfileģ������
	regfile regfile1(
		.clk(clk),
		.rst(rst),
		.we(wb_wreg_i),
		.waddr(wb_wd_i),
		.wdata(wb_wdata_i),
		.re1(reg1_read),
		.raddr1(reg1_addr),
		.rdata1(reg1_data),
		.re2(reg2_read),
		.raddr2(reg2_addr),
		.rdata2(reg2_data),
		.select(select[4:0]),
		.output_data(regfile_data_o)
	);

	//ID/EXģ������
	id_ex id_ex0(
		.clk(clk),
		.rst(rst),

		.stall(stall),
		.flush(flush),

		//������׶�IDģ�鴫�ݹ�������Ϣ
		.id_aluop(id_aluop_o),
		.id_alusel(id_alusel_o),
		.id_reg1(id_reg1_o),
		.id_reg2(id_reg2_o),
		.id_wd(id_wd_o),
		.id_wreg(id_wreg_o),
		.id_link_address(id_link_address_o),
		.id_is_in_delayslot(id_is_in_delayslot_o),
		.next_inst_in_delayslot_i(next_inst_in_delayslot_o),
		.id_inst(id_inst_o),
		.id_excepttype(id_excepttype_o),
		.id_current_inst_address(id_current_inst_address_o),

		//���ݵ�ִ�н׶�EXģ�����Ϣ
		.ex_aluop(ex_aluop_i),
		.ex_alusel(ex_alusel_i),
		.ex_reg1(ex_reg1_i),
		.ex_reg2(ex_reg2_i),
		.ex_wd(ex_wd_i),
		.ex_wreg(ex_wreg_i),
		.ex_link_address(ex_link_address_i),
		.ex_is_in_delayslot(ex_is_in_delayslot_i),
		.is_in_delayslot_o(is_in_delayslot_i),
		.ex_inst(ex_inst_i),
		.ex_excepttype(ex_excepttype_i),
		.ex_current_inst_address(ex_current_inst_address_i)
	);

	//EXģ������
	ex ex0(
		.rst(rst),

		//��ID/EXģ�鴫�ݹ�������Ϣ
		.aluop_i(ex_aluop_i),
		.alusel_i(ex_alusel_i),
		.reg1_i(ex_reg1_i),
		.reg2_i(ex_reg2_i),
		.wd_i(ex_wd_i),
		.wreg_i(ex_wreg_i),
		.hi_i(hi),
		.lo_i(lo),
		.inst_i(ex_inst_i),

		//�����EX/MEMģ�����Ϣ
		.wb_hi_i(wb_hi_i),
		.wb_lo_i(wb_lo_i),
		.wb_whilo_i(wb_whilo_i),
		.mem_hi_i(mem_hi_o),
		.mem_lo_i(mem_lo_o),
		.mem_whilo_i(mem_whilo_o),

		.link_address_i(ex_link_address_i),
		.is_in_delayslot_i(ex_is_in_delayslot_i),

		.excepttype_i(ex_excepttype_i),
		.current_inst_address_i(ex_current_inst_address_i),

		//�ô�׶ε�ָ���Ƿ�ҪдCP0����������������
		.mem_cp0_reg_we(mem_cp0_reg_we_o),
		.mem_cp0_reg_write_addr(mem_cp0_reg_write_addr_o),
		.mem_cp0_reg_data(mem_cp0_reg_data_o),

		//��д�׶ε�ָ���Ƿ�ҪдCP0����������������
		.wb_cp0_reg_we(wb_cp0_reg_we_i),
		.wb_cp0_reg_write_addr(wb_cp0_reg_write_addr_i),
		.wb_cp0_reg_data(wb_cp0_reg_data_i),

		.cp0_reg_data_i(cp0_data_o),
		.cp0_reg_read_addr_o(cp0_raddr_i),
		
		//����һ��ˮ�����ݣ�����дCP0�еļĴ���
		.cp0_reg_we_o(ex_cp0_reg_we_o),
		.cp0_reg_write_addr_o(ex_cp0_reg_write_addr_o),
		.cp0_reg_data_o(ex_cp0_reg_data_o),

		.wd_o(ex_wd_o),
		.wreg_o(ex_wreg_o),
		.wdata_o(ex_wdata_o),
		.hi_o(ex_hi_o),
		.lo_o(ex_lo_o),
		.whilo_o(ex_whilo_o),

		.aluop_o(ex_aluop_o),
		.mem_addr_o(ex_mem_addr_o),
		.reg2_o(ex_reg2_o),
		
		.excepttype_o(ex_excepttype_o),
		.is_in_delayslot_o(ex_is_in_delayslot_o),
		.current_inst_address_o(ex_current_inst_address_o),
		.stallreq(stallreq_from_ex)
	);

	//EX/MEMģ������
	ex_mem ex_mem0(
		.clk(clk),
		.rst(rst),
		.stall(stall),
		.flush(flush),

		//����ִ�н׶�EXģ�����Ϣ
		.ex_wd(ex_wd_o),
		.ex_wreg(ex_wreg_o),
		.ex_wdata(ex_wdata_o),
		.ex_hi(ex_hi_o),
		.ex_lo(ex_lo_o),
		.ex_whilo(ex_whilo_o),

		.ex_aluop(ex_aluop_o),
		.ex_mem_addr(ex_mem_addr_o),
		.ex_reg2(ex_reg2_o),

		.ex_cp0_reg_we(ex_cp0_reg_we_o),
		.ex_cp0_reg_write_addr(ex_cp0_reg_write_addr_o),
		.ex_cp0_reg_data(ex_cp0_reg_data_o),

		.ex_excepttype(ex_excepttype_o),
		.ex_is_in_delayslot(ex_is_in_delayslot_o),
		.ex_current_inst_address(ex_current_inst_address_o),

		//�͵��ô�׶�MEMģ�����Ϣ
		.mem_wd(mem_wd_i),
		.mem_wreg(mem_wreg_i),
		.mem_wdata(mem_wdata_i),
		.mem_hi(mem_hi_i),
		.mem_lo(mem_lo_i),
		.mem_whilo(mem_whilo_i),

		.mem_cp0_reg_we(mem_cp0_reg_we_i),
		.mem_cp0_reg_write_addr(mem_cp0_reg_write_addr_i),
		.mem_cp0_reg_data(mem_cp0_reg_data_i),

		.mem_aluop(mem_aluop_i),
		.mem_mem_addr(mem_mem_addr_i),
		.mem_reg2(mem_reg2_i),

		.mem_excepttype(mem_excepttype_i),
		.mem_is_in_delayslot(mem_is_in_delayslot_i),
		.mem_current_inst_address(mem_current_inst_address_i)
	);

	//MEMģ������
	mem mem0(
		.rst(rst),

		//����EX/MEMģ�����Ϣ
		.wd_i(mem_wd_i),
		.wreg_i(mem_wreg_i),
		.wdata_i(mem_wdata_i),
		.hi_i(mem_hi_i),
		.lo_i(mem_lo_i),
		.whilo_i(mem_whilo_i),

		.aluop_i(mem_aluop_i),
		.mem_addr_i(mem_mem_addr_i),
		.reg2_i(mem_reg2_i),

		.mem_data_i(ram_data_i),

		.cp0_reg_we_i(mem_cp0_reg_we_i),
		.cp0_reg_write_addr_i(mem_cp0_reg_write_addr_i),
		.cp0_reg_data_i(mem_cp0_reg_data_i),

		.excepttype_i(mem_excepttype_i),
		.is_in_delayslot_i(mem_is_in_delayslot_i),
		.current_inst_address_i(mem_current_inst_address_i),

		.cp0_bad_v_addr_i(cp0_bad_v_addr),
		.cp0_status_i(cp0_status),
		.cp0_cause_i(cp0_cause),
		.cp0_epc_i(cp0_epc),
		.cp0_index_i(cp0_index),
		.cp0_entry_lo_0_i(cp0_entry_lo_0),
		.cp0_entry_lo_1_i(cp0_entry_lo_1),
		.cp0_entry_hi_i(cp0_entry_hi),

		//��д�׶ε�ָ���Ƿ�ҪдCP0����������������
		.wb_cp0_reg_we(wb_cp0_reg_we_i),
		.wb_cp0_reg_write_addr(wb_cp0_reg_write_addr_i),
		.wb_cp0_reg_data(wb_cp0_reg_data_i),

		.excepttype_is_tlbm_i(tlb_excepttype_is_tlbm),
		.excepttype_is_tlbl_i(tlb_excepttype_is_tlbl),
		.excepttype_is_tlbs_i(tlb_excepttype_is_tlbs),

		//�͵�CP0ģ�����Ϣ
		.cp0_reg_we_o(mem_cp0_reg_we_o),
		.cp0_reg_write_addr_o(mem_cp0_reg_write_addr_o),
		.cp0_reg_data_o(mem_cp0_reg_data_o),

		.excepttype_o(mem_excepttype_o),
		.cp0_epc_o(latest_epc),
		.is_in_delayslot_o(mem_is_in_delayslot_o),
		.current_inst_address_o(mem_current_inst_address_o),
		.bad_v_addr_o(bad_v_addr_o),

		//�͵�MEM/WBģ�����Ϣ
		.wd_o(mem_wd_o),
		.wreg_o(mem_wreg_o),
		.wdata_o(mem_wdata_o),
		.hi_o(mem_hi_o),
		.lo_o(mem_lo_o),
		.whilo_o(mem_whilo_o),

		//�͵�MMUģ�����Ϣ
		.mem_addr_o(ram_addr_o),
		.mem_we_o(ram_we_o),
		.mem_sel_o(ram_sel_o),
		.mem_data_o(ram_data_o),
		.mem_ce_o(ram_ce_o),

		//�͵�TLBģ�����Ϣ
		.tlb_we_o(tlb_we),
		.tlb_index_o(tlb_index),
		.tlb_data_o(tlb_data)
	);

	//MEM/WBģ������
	mem_wb mem_wb0(
		.clk(clk),
		.rst(rst),
		.stall(stall),
		.flush(flush),
		
		//���Էô�׶�MEMģ�����Ϣ
		.mem_wd(mem_wd_o),
		.mem_wreg(mem_wreg_o),
		.mem_wdata(mem_wdata_o),
		.mem_hi(mem_hi_o),
		.mem_lo(mem_lo_o),
		.mem_whilo(mem_whilo_o),

		.mem_cp0_reg_we(mem_cp0_reg_we_o),
		.mem_cp0_reg_write_addr(mem_cp0_reg_write_addr_o),
		.mem_cp0_reg_data(mem_cp0_reg_data_o),

		//�͵���д�׶ε���Ϣ
		.wb_wd(wb_wd_i),
		.wb_wreg(wb_wreg_i),
		.wb_wdata(wb_wdata_i),
		.wb_hi(wb_hi_i),
		.wb_lo(wb_lo_i),
		.wb_whilo(wb_whilo_i),
		
		.wb_cp0_reg_we(wb_cp0_reg_we_i),
		.wb_cp0_reg_write_addr(wb_cp0_reg_write_addr_i),
		.wb_cp0_reg_data(wb_cp0_reg_data_i)
	);

	hilo_reg hilo_reg0(
		.clk(clk),
		.rst(rst),

		//д�˿�
		.we(wb_whilo_i),
		.hi_i(wb_hi_i),
		.lo_i(wb_lo_i),

		//���˿�1
		.hi_o(hi),
		.lo_o(lo)
	);

	ctrl ctrl0(
		.rst(rst),

		.excepttype_i(mem_excepttype_o),
		.cp0_epc_i(latest_epc),
	
		.stallreq_from_if(stallreq_from_if),
		.stallreq_from_id(stallreq_from_id),
		.stallreq_from_ex(stallreq_from_ex),
		.stallreq_from_mem(stallreq_from_mem),

		.new_pc(new_pc),
		.flush(flush),
		.stall(stall)
	);

	cp0_reg cp0_reg0(
		.clk(clk),
		.rst(rst),

		.we_i(wb_cp0_reg_we_i),
		.waddr_i(wb_cp0_reg_write_addr_i),
		.raddr_i(cp0_raddr_i),
		.data_i(wb_cp0_reg_data_i),

		.excepttype_i(mem_excepttype_o),
		.int_i(int_i),
		.current_inst_addr_i(mem_current_inst_address_o),
		.bad_v_addr_i(bad_v_addr_o),
		.is_in_delayslot_i(mem_is_in_delayslot_o),

		.data_o(cp0_data_o),
		.index_o(cp0_index),
		.entry_lo_0_o(cp0_entry_lo_0),
		.entry_lo_1_o(cp0_entry_lo_1),
		.bad_v_addr_o(cp0_bad_v_addr),
		.count_o(cp0_count),
		.entry_hi_o(cp0_entry_hi),
		.compare_o(cp0_compare),
		.status_o(cp0_status),
		.cause_o(cp0_cause),
		.epc_o(cp0_epc),
		.ebase_o(cp0_ebase),
		
		.timer_int_o(timer_int_o)
	);

	mmu mmu0(
		.clk(clk),
		.rst(rst),

		.tlb_addr_i(tlb_addr_i),

		.mmu_addr_o(mmu_addr_i),
		.mmu_select_o(mmu_select_i)
	);

	tlb tlb0(
		.clk(clk),
		.rst(rst),

		.bus_addr_i(bus_addr_i),
		.bus_write_i(bus_write_i),
		.tlb_ce(tlb_ce_i),
		.tlb_addr(tlb_addr_i),

		.tlb_we(tlb_we),
		.tlb_index(tlb_index),
		.tlb_data(tlb_data),

		.excepttype_is_tlbm(tlb_excepttype_is_tlbm),
		.excepttype_is_tlbl(tlb_excepttype_is_tlbl),
		.excepttype_is_tlbs(tlb_excepttype_is_tlbs)
	);

	wishbone_bus wishbone_bus0(
		.clk(clk),
		.rst(rst),

		//���Կ���ģ��Ctrl
		.stall_i(stall),
		.flush_i(flush),

		//IFģ��Ľӿ�
		.if_ce_i(rom_ce),
		.if_data_i(32'h00000000),
		.if_addr_i(next_pc),
		.if_we_i(1'b0),
		.if_sel_i(4'b1111),
		.if_data_o(inst_i),

		.stall_req_if(stallreq_from_if),

		//MEMģ��Ľӿ�
		.mem_ce_i(ram_ce_o),
		.mem_data_i(ram_data_o),
		.mem_addr_i(ram_addr_o),
		.mem_we_i(ram_we_o),
		.mem_sel_i(ram_sel_o),
		.mem_data_o(ram_data_i),

		.stall_req_mem(stallreq_from_mem),

		//TLBģ��Ľӿ�
		.tlb_write_o(bus_write_i),
		.tlb_ce(tlb_ce_i),
		.tlb_addr_o(bus_addr_i),

		//MMUģ��Ľӿ�
		.mmu_addr_i(mmu_addr_i),
		.mmu_select_i(mmu_select_i),

		//Wishbone���߲�ӿ�
		.wishbone_data_i(wishbone_data_i),
		.wishbone_ack_i(wishbone_ack_i),
		.wishbone_addr_o(wishbone_addr_o),
		.wishbone_data_o(wishbone_data_o),
		.wishbone_we_o(wishbone_we_o),
		.wishbone_select_o(wishbone_select_o),
		.state(state)
	);

endmodule
